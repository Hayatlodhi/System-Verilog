int arr[3] = '{5,6,7};  // Declaration, and assignment
Or
int arr[3];
arr[0] = 5;
arr[1] = 6;
arr[2] = 7;

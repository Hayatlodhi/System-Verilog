// declaration of array 
int arr[2] = '{3,4};  // Declaration, and assignment
Or
int arr[2];
arr[0] = 3;
arr[1] = 4;
